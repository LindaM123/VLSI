**.subckt sim_inv1
x1 vdd vin vout vss inv1
C1 vout GND 10f m=1
V1 vin GND PULSE(0 1.8 2n 10p 10p 2n 4n)
V2 vdd GND 1.8
V3 vss GND 0
**** begin user architecture code



.lib ~/tecnicas_digitales_programas/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.control
set color0 = rgb:f/f/e
tran 0.01ns 5n
plot vin vout
.endc

.save all



**** end user architecture code
**.ends

* expanding   symbol:  inv1.sym # of pins=4
* sym_path: /home/julious/tecnicas_digitales_programas/inversor_simulacion/inv1.sym
* sch_path: /home/julious/tecnicas_digitales_programas/inversor_simulacion/inv1.sch
.subckt inv1  Vdd! in out Vss!
*.iopin Vdd!
*.iopin Vss!
*.ipin in
*.opin out
XM1 out in Vss! Vss! sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 out in Vdd! Vdd! sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

.GLOBAL GND
** flattened .save nodes
.end
